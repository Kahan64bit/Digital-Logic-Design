//NOT gate using Structural modeling
module not_gate_s(a,y);
 input a;
 output y;

 not(y,a);

endmodule